module shifter (A, B, SL, SR);

input [31:0] A, B;

output [31:0] SL, SR;


endmodule
